library verilog;
use verilog.vl_types.all;
entity Clock_Devider_vlg_check_tst is
    port(
        CLK_1ms         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Clock_Devider_vlg_check_tst;
