library verilog;
use verilog.vl_types.all;
entity Clock_Devider_vlg_vec_tst is
end Clock_Devider_vlg_vec_tst;
