library verilog;
use verilog.vl_types.all;
entity System_vlg_vec_tst is
end System_vlg_vec_tst;
