library verilog;
use verilog.vl_types.all;
entity Led_Control_vlg_vec_tst is
end Led_Control_vlg_vec_tst;
