library verilog;
use verilog.vl_types.all;
entity Clock_Devider_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Clock_Devider_vlg_sample_tst;
